lmao = ptdr