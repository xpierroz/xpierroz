wouaf = bruh
xxx = test
jklm = xxf