AutoRep DM | 3/09/21 - 16:43:30 - .$ - 765850375965638686 - .$'s server - 808250457847234570 - lmao - ptdrAutoRep DM | 3/09/21 - 17:30:10 - .$ - 765850375965638686 - .$'s server - 808250457847234570 - lmao - ptdrAutoRep DM | 3/11/21 - 15:42:51 - .$ - 819487357904355360 - .$'s server - 808250457847234570 - lmao - ptdr
AutoRep DM | 03/11/21 13:53:11 - .$ - 819487357904355360 - .$'s server - 808250457847234570 - lmao - ptdr
